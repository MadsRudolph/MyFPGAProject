----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:32:05 05/05/2025 
-- Design Name: 
-- Module Name:    Sawtooth - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEE.STD_LOGIC_unsigned.ALL;

entity Sawtooth is
    Port ( Reset : in  STD_LOGIC;
           Clk : in  STD_LOGIC;
           SigAmpl : out  STD_LOGIC);
end Sawtooth;

architecture Behavioral of Sawtooth is

begin

Sawtooth: process()

end Behavioral;

